-- http://jacques.weber.pagesperso-orange.fr/vhdl_html/Vhdl.htm
-- http://hdl.telecom-paristech.fr/vhdl_structurel.html
-- http://amouf.chez.com/syntaxe.htm

library IEEE;	-- type boolean, bit, character, severity_level
use IEEE.STD_LOGIC_1164.ALL;	-- definit les types std_logic , std_logic_vector , std_ulogic, les opérateurs logiques et les fonctions de recherches de fronts rising_edge() et falling_edge(). introduit par IEE 1164 en 1992.
use IEEE.NUMERIC_STD.ALL;		-- definit les sous-types entier "signed" ou "unsigned", introduit par IEEE 1076.3
use IEEE.NUMERIC_BIT.ALL; 		-- définit les opérateurs arithmétiques agissant sur des bit_vector interprétés comme des nombres entiers.
use std.textio.all; 
use IEEE.std_logic_arith, IEEE.std_logic_misc, IEEE.std_logic_signed, IEEE.std_logic_textio, IEEE.std_logic_unsigned -- ancienne librairie par IEEE de 1989.

Constant T_PD : time := 5 ns ;

entity nom_entity is
-- generic (n: natural:=32);		
port( 					-- (rappel: le dernier listing de port n'a pas de ;)
		a,b : in unsigned(2 downto 0);  
        c : out std_logic; 
        d : in std_logic;  
        a_gt_b : out std_logic  
      );    
end nom_entity;

architecture nom_archi of nom_entity is

-- example declatation signal avec valeur par default: signal temp1,temp2,temp3 : std_logic := '0';
-- example declaration signal avec range: signal i : integer range 0 to 30:=0;
type memory_type is array (0 to 29) of integer range -128 to 127;
--ROM for storing the sine values generated by MATLAB.
signal sine : memory_type :=(0,16,31,45,58,67,74,77,77,74,67,58,45,31,16,0,
-16,-31,-45,-58,-67,-74,-77,-77,-74,-67,-58,-45,-31,-16);

BEGIN

-- example affectation:	temp1 <= not(a(2) xor b(2));  --XNOR gate with 2 inputs.
-- example affectation tableau1: temp(1) <= temp(0);
-- example affectation tableau2: temp <= (0=> '1', others => '0');
-- example décalage: a:=adecaler ror decombien; b:=adecaler rol decombien;
-- opérateurs logiques:  and | or | nand | nor | xor | xnor
-- Opérateurs relationnels:  = | /= | < | <= | > | >=
-- Opérateurs de décalage: sll | srl | sla | sra | rol | ror
-- Opérateurs d’addition:  + | – | 
-- operateur de concaténation: &
-- Opérateurs de multiplication: * | / | mod | rem
-- 		mod : quotient division euclidienne
--		rem : reste division euclidienne     A = (A mod b) * b + (a rem b)
-- Opérateurs divers:  ** | abs | not

process(CLR,PRE,CLK) --process with sensitivity list.
begin  --"begin" statment for the process.

-- if
    if (CLR = '1') then  --Asynchronous clear input
           Q <= '0';
    else
           if(PRE = '1') then  --Asynchronous set input
               Q <= '1';
           else
               if ( CE = '1' and  falling_edge(CLK) ) then
                  Q <= D;      
              end if;
          end if;
   end if;
   
if condition1 then
--- instructions séquentielles 1
[elsif condition2 then
--- instructions séquentielles 2]
[elsif condition3 then
--- instructions séquentielles 3]
[else
--- instructions séquentielles n]
end if ;

-- boucle while   *** Attention: la boucle while n'est pas synthetisable
While condition Loop
		listeInstructionsSéquentielles
end loop ;

-- boucle for
for identifiantVariable in gammeDiscrète loop
		listeInstructionsSéquentielles
end loop ; 

-- boucle case
case expression is
	when choix =>
		listeInstructionsSéquentielles
	…
	when choix =>
		listeInstructionsSéquentielles
	when others =>
		listeInstructionsSéquentielles
end case;

-- with select
with cmd select
	q <= 	bus0 when "00",
			bus1 when "01",
			bus2 when "10",
			bus3 when "11",
			bus0 when others;

end process;  --end of process statement.

end nom_archi;